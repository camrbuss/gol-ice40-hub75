// MIT License

// Copyright (c) [2021] [camrbuss]

// Permission is hereby granted, free of charge, to any person obtaining a copy
// of this software and associated documentation files (the "Software"), to deal
// in the Software without restriction, including without limitation the rights
// to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
// copies of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:

// The above copyright notice and this permission notice shall be included in all
// copies or substantial portions of the Software.

// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
// IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
// FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
// AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
// LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
// OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
// SOFTWARE.


// To use the test bench with iverilog you will need to switch the 24 mHz clock
// to a clk generated by the test bench as the simulation of the pll does not
// generate a clock. Other than the clock there are no other inputs.

module top
(
    // input clk,
	output reg R0,
	output reg G0,
	output reg B0,
	output reg B1,
	output reg G1,
	output reg R1,
	output reg A0,
	output reg A1,
	output reg A2,
	output reg A3,
	output reg A4,
	output reg CK,
	output reg LA,
	output reg BL);

reg [15:0] P_DAT0 [255:0];
reg [15:0] P_DAT1 [255:0];
reg [15:0] P_DAT2 [255:0];
reg [15:0] P_DAT3 [255:0];
reg [15:0] P_DAT4 [255:0];
reg [15:0] P_DAT5 [255:0];
reg [15:0] P_DAT6 [255:0];
reg [15:0] P_DAT7 [255:0];

// Initialize the plls for 24 mHz clocked output to the matrix
wire clk_48mhz;
wire clk_24mhz;
SB_HFOSC SB_HFOSC_inst(
	.CLKHFEN(1'b1),
	.CLKHFPU(1'b1),
	.CLKHF(clk_48mhz)
);
SB_PLL40_CORE #(
	.FEEDBACK_PATH("SIMPLE"),
	.PLLOUT_SELECT("GENCLK"),
	.DIVR(4'b0000),
	.DIVF(7'b0001111),
	.DIVQ(3'b101),
	.FILTER_RANGE(3'b100)
) SB_PLL40_CORE_inst (
	.RESETB(1'b1),
	.BYPASS(1'b0),
	.PLLOUTCORE(clk_24mhz),
	.REFERENCECLK(clk_48mhz)
);

// os = ongoing state
// os_t = ongoing state top (first 32 rows)
// os_b = ongoing state bot (bottom 32 rows)
// each address contains 1/4 of a row
// Address  0                1                2                3
// Data     1111111111111111 1111111111111111 1111111111111111 1111111111111111
// Address  4                5                6                7
// Data     1111111111111111 1111111111111111 1111111111111111 1111111111111111
//          ... all the way to address 255

// ns_spram = next state
// Each address only holds data in the first bit position.
// This way the address can be used to get the neighboring cells
// of the current cell that is being evaluated

reg [13:0] os_addr = 0;
reg [13:0] os_disp_addr;
reg [13:0] os_gol_addr;
reg [15:0] os_t_data_in = 0;
reg [15:0] os_b_data_in = 0;
reg os_t_wren;
reg os_b_wren;
wire [15:0] os_t_data_out;
wire [15:0] os_b_data_out;

reg [11:0] ns_addr = 0;
reg [15:0] ns_data_in;
reg ns_wren = 0;
wire [15:0] ns_data_out;

SB_SPRAM256KA os_t_spram
(
	.ADDRESS(os_addr),
	.DATAIN(os_t_data_in),
	.MASKWREN({os_t_wren, os_t_wren, os_t_wren, os_t_wren}),
	.WREN(os_t_wren),
	.CHIPSELECT(1'b1),
	.CLOCK(clk_24mhz),
	.STANDBY(1'b0),
	.SLEEP(1'b0),
	.POWEROFF(1'b1),
	.DATAOUT(os_t_data_out)
);

SB_SPRAM256KA os_b_spram
(
	.ADDRESS(os_addr),
	.DATAIN(os_b_data_in),
	.MASKWREN({os_b_wren, os_b_wren, os_b_wren, os_b_wren}),
	.WREN(os_b_wren),
	.CHIPSELECT(1'b1),
	.CLOCK(clk_24mhz),
	.STANDBY(1'b0),
	.SLEEP(1'b0),
	.POWEROFF(1'b1),
	.DATAOUT(os_b_data_out)
);

SB_SPRAM256KA ns_spram
(
	.ADDRESS(ns_addr),
	.DATAIN(ns_data_in),
	.MASKWREN({ns_wren, ns_wren, ns_wren, ns_wren}),
	.WREN(ns_wren),
	.CHIPSELECT(1'b1),
	.CLOCK(clk_24mhz),
	.STANDBY(1'b0),
	.SLEEP(1'b0),
	.POWEROFF(1'b1),
	.DATAOUT(ns_data_out)
);

reg [6:0] preload_cnt = 0;
reg [2:0] preload_switch = 0;
reg [15:0] tcol0;
reg [15:0] tcol1;
reg [15:0] tcol2;
reg [15:0] tcol3;
reg [15:0] bcol0;
reg [15:0] bcol1;
reg [15:0] bcol2;
reg [15:0] bcol3;

reg [11:0] idx = 0;  // 64 * 64 = 4096 positions
reg [3:0] population = 0;
reg curr_state = 0;
reg [31:0] gol_state = 0;
reg [13:0] cycles = 0;
reg [3:0] neigh = 4'b1111;
reg [11:0] neigh_addr;
reg [15:0] block_buff;

// TODO: convert numbers to enumerations?
always @(posedge clk_24mhz) begin
	case (gol_state)
		0: begin
			os_addr <= preload_cnt;
			case (preload_switch)
				3'b000: begin
					os_t_data_in <= P_DAT0[preload_cnt];
					os_b_data_in <= P_DAT0[preload_cnt+128];
				end
				3'b001: begin
					os_t_data_in <= P_DAT1[preload_cnt];
					os_b_data_in <= P_DAT1[preload_cnt+128];
				end
				3'b010: begin
					os_t_data_in <= P_DAT2[preload_cnt];
					os_b_data_in <= P_DAT2[preload_cnt+128];
				end
				3'b011: begin
					os_t_data_in <= P_DAT3[preload_cnt];
					os_b_data_in <= P_DAT3[preload_cnt+128];
				end
				3'b100: begin
					os_t_data_in <= P_DAT4[preload_cnt];
					os_b_data_in <= P_DAT4[preload_cnt+128];
				end
				3'b101: begin
					os_t_data_in <= P_DAT5[preload_cnt];
					os_b_data_in <= P_DAT5[preload_cnt+128];
				end
				3'b110: begin
					os_t_data_in <= P_DAT6[preload_cnt];
					os_b_data_in <= P_DAT6[preload_cnt+128];
				end
				3'b111: begin
					os_t_data_in <= P_DAT7[preload_cnt];
					os_b_data_in <= P_DAT7[preload_cnt+128];
				end
				default: begin
					os_t_data_in <= P_DAT0[preload_cnt];
					os_b_data_in <= P_DAT0[preload_cnt+128];
				end
			endcase

			os_t_wren <= 1;
			os_b_wren <= 1;
			preload_cnt <= preload_cnt + 1;
			if (preload_cnt == 7'b1111111) begin
				gol_state <= gol_state + 1;
			end
		end
		1: begin
			os_t_wren <= 0;
			os_b_wren <= 0;
			os_addr <= idx[10:4];
			gol_state <= gol_state + 1;
		end
		2: begin
			gol_state <= gol_state + 1;
		end
		3: begin
			gol_state <= gol_state + 1;
		end
		4: begin
			ns_wren <= 1;
			ns_addr <= idx;
			if (idx[11] == 0) begin
				ns_data_in <= os_t_data_out[15-idx[3:0]];
			end else begin
				ns_data_in <= os_b_data_out[15-idx[3:0]];
			end
			idx <= idx + 1;
			if (idx == 12'b111111111111) begin
				gol_state <= gol_state + 1;
			end else if (idx[3:0] == 4'b1111) begin
				gol_state <= 1;
			end
		end
		5: begin
			ns_wren <= 0;
			gol_state <= gol_state + 1;
			idx <= 0;
		end
		6: begin
			gol_state <= gol_state + 1;
			neigh <= 4'b1111;
		end
		7: begin
			os_t_wren <= 0;
			os_b_wren <= 0;
			case (neigh)
				0: ns_addr <= idx;
				1: ns_addr <= idx - 65; // Top left
				2: ns_addr <= idx - 64; // Top
				3: ns_addr <= idx - 63; // Top Right
				4: ns_addr <= idx - 1; // Left
				5: ns_addr <= idx + 1; // Right
				6: ns_addr <= idx + 65; // Bot Right
				7: ns_addr <= idx + 64; // Bot
				8: ns_addr <= idx + 63; // Bot Left
				default: begin
					// gol_state <= 5;
					neigh <= 8;
					population <= 0;
					idx <= idx + 1;
				end
			endcase
			if (neigh > 8) begin
				gol_state <= 7;
			end else begin
				gol_state <= gol_state + 1;
			end
		end
		8: begin
			if (ns_addr > 4095) begin
				if (neigh < 5) begin
					ns_addr <= 4096 - (4096 - neigh);
				end else begin
					ns_addr <= ns_addr - 4096;
				end
			end else begin
				gol_state <= gol_state + 1;
			end
		end
		9: begin
			gol_state <= gol_state + 1;
		end
		10: begin
			if (neigh == 0) begin
				// Determine if the cell should live or die
				if (population == 3 || (population == 2 && ns_data_out[0] == 1)) begin
					block_buff[15-idx[3:0]] <= 1'b1;
				end else begin
					block_buff[15-idx[3:0]] <= 1'b0;
				end
			end else begin
				population <= population + ns_data_out[0];
			end

			if (idx[3:0] == 4'b1111 && neigh[3:0] == 4'b0000) begin
				// push the block_buff into displayed spram
				gol_state <= gol_state + 1;
				os_addr <= idx[10:4];
			end else begin
				gol_state <= 7;
			end
			neigh <= neigh - 1;
		end
		11: begin
			gol_state <= gol_state + 1;
		end
		12: begin
			if (idx[11] == 0) begin
				os_t_wren <= 1;
				os_t_data_in <= block_buff;
			end else begin
				os_b_wren <= 1;
				os_b_data_in <= block_buff;
			end
			gol_state <= gol_state + 1;
		end
		13: begin
			os_t_wren <= 0;
			os_b_wren <= 0;
			os_addr <= os_addr + 1;
			if (idx == 12'b111111111111) begin
				// gol_state <= 0;
				gol_state <= gol_state + 1;
				idx <= 0;
			end else begin
				gol_state <= 7;
			end
		end
		// The value of this case determines the play rate
		// 32'hFFFFFFFF: begin
		32'h000FFFFF: begin
		// 100: begin
			gol_state <= 1;
            cycles <= cycles + 1;
			// The number of bits from cycles determines the rate at which
			// the preload value changes
            if (preload_switch != cycles[13:11]) begin
				preload_switch <= cycles[13:11];
				gol_state <= 0;
			end
		end

		default: begin
			gol_state <= gol_state + 1;
			os_t_wren <= 0;
			os_b_wren <= 0;
			os_addr <= os_disp_addr;

		end
	endcase

end


reg [63:0] r0 = 0;
reg [63:0] r1 = 0;
reg [15:0] r0_c0 = 0;
reg [15:0] r0_c1 = 0;
reg [15:0] r0_c2 = 0;
reg [15:0] r0_c3 = 0;
reg [15:0] r1_c0 = 0;
reg [15:0] r1_c1 = 0;
reg [15:0] r1_c2 = 0;
reg [15:0] r1_c3 = 0;

reg [4:0] address = 0; // Vertical Address
reg [6:0] state = 0;
reg half_div = 0;
reg [5:0] horiz_cnt = 0; // Horizontal "Address"

initial begin

	R0         = 0;
	G0         = 0;
	B0         = 0;
	B1         = 0;
	G1         = 0;
	R1         = 0;
	LA         = 0;
	BL         = 0;
	A0         = 0; // LSB
	A1         = 0;
	A2         = 0;
	A3         = 0;
	A4         = 0; // MSB
	CK         = 0;

	// Randomn MWSS's
	P_DAT0[0] = 16'b1111000000000000; P_DAT0[1] = 16'b0000000000000000; P_DAT0[2] = 16'b0000000000000000; P_DAT0[3] = 16'b0000000000000000;
	P_DAT0[4] = 16'b0000000000000000; P_DAT0[5] = 16'b0000000000000000; P_DAT0[6] = 16'b0000000000000000; P_DAT0[7] = 16'b0000000000000000;
	P_DAT0[8] = 16'b0000000000000000; P_DAT0[9] = 16'b0000000000000000; P_DAT0[10] = 16'b0000000000000000; P_DAT0[11] = 16'b0000000000000000;
	P_DAT0[12] = 16'b0000110000000000; P_DAT0[13] = 16'b0001111000000000; P_DAT0[14] = 16'b0000110000000000; P_DAT0[15] = 16'b0000110000000000;
	P_DAT0[16] = 16'b0001101110000000; P_DAT0[17] = 16'b0001111110000000; P_DAT0[18] = 16'b0001101110000000; P_DAT0[19] = 16'b0001101110000000;
	P_DAT0[20] = 16'b0000111110000000; P_DAT0[21] = 16'b0000111110000000; P_DAT0[22] = 16'b0000111110000000; P_DAT0[23] = 16'b0000111110000000;
	P_DAT0[24] = 16'b0000011100000000; P_DAT0[25] = 16'b0000011100000000; P_DAT0[26] = 16'b0000011100000000; P_DAT0[27] = 16'b0000011100000000;
	P_DAT0[28] = 16'b0000000000000000; P_DAT0[29] = 16'b0000000000000000; P_DAT0[30] = 16'b0000000000000000; P_DAT0[31] = 16'b0000000000000000;
	P_DAT0[32] = 16'b0000000000000000; P_DAT0[33] = 16'b0000000000000000; P_DAT0[34] = 16'b0000000000000000; P_DAT0[35] = 16'b0000000000000000;
	P_DAT0[36] = 16'b0000000000000000; P_DAT0[37] = 16'b0000000000000000; P_DAT0[38] = 16'b0000000000000000; P_DAT0[39] = 16'b0000010100000000;
	P_DAT0[40] = 16'b0000111000000000; P_DAT0[41] = 16'b0000000000000000; P_DAT0[42] = 16'b0000000000000000; P_DAT0[43] = 16'b0000001000000000;
	P_DAT0[44] = 16'b0000111000000000; P_DAT0[45] = 16'b0000000000000000; P_DAT0[46] = 16'b0000000000000000; P_DAT0[47] = 16'b0000010100000000;
	P_DAT0[48] = 16'b0000111000000000; P_DAT0[49] = 16'b0000000000000000; P_DAT0[50] = 16'b0000000000000000; P_DAT0[51] = 16'b0000000000000000;
	P_DAT0[52] = 16'b0000000000000000; P_DAT0[53] = 16'b0000000000000000; P_DAT0[54] = 16'b0000000000000000; P_DAT0[55] = 16'b0000000000000000;
	P_DAT0[56] = 16'b0000000000000000; P_DAT0[57] = 16'b0000000000000000; P_DAT0[58] = 16'b0000000000000000; P_DAT0[59] = 16'b0000000000000000;
	P_DAT0[60] = 16'b0000000000000000; P_DAT0[61] = 16'b0000000000000000; P_DAT0[62] = 16'b0000000000000000; P_DAT0[63] = 16'b0000000000000000;
	P_DAT0[64] = 16'b0000000000000000; P_DAT0[65] = 16'b0000000000000000; P_DAT0[66] = 16'b0000000000000000; P_DAT0[67] = 16'b0000000000000000;
	P_DAT0[68] = 16'b0000000000000000; P_DAT0[69] = 16'b0000000000000000; P_DAT0[70] = 16'b0000000000000000; P_DAT0[71] = 16'b0000000000000000;
	P_DAT0[72] = 16'b0000000000000000; P_DAT0[73] = 16'b0000000000000000; P_DAT0[74] = 16'b0000000000000000; P_DAT0[75] = 16'b0000000000000000;
	P_DAT0[76] = 16'b0000110000000000; P_DAT0[77] = 16'b0000110000000000; P_DAT0[78] = 16'b0000110000000000; P_DAT0[79] = 16'b0000110000000000;
	P_DAT0[80] = 16'b0001101110000000; P_DAT0[81] = 16'b0001101110000000; P_DAT0[82] = 16'b0001101110000000; P_DAT0[83] = 16'b0001101110000000;
	P_DAT0[84] = 16'b0000111110000000; P_DAT0[85] = 16'b0000111110000000; P_DAT0[86] = 16'b0000111110000000; P_DAT0[87] = 16'b0000111110000000;
	P_DAT0[88] = 16'b0000011100000000; P_DAT0[89] = 16'b0000011100000000; P_DAT0[90] = 16'b0000011100000000; P_DAT0[91] = 16'b0000011100000000;
	P_DAT0[92] = 16'b0000000000000000; P_DAT0[93] = 16'b0000000000000000; P_DAT0[94] = 16'b0000000000000000; P_DAT0[95] = 16'b0000000000000000;
	P_DAT0[96] = 16'b0000000000000000; P_DAT0[97] = 16'b0000000000000000; P_DAT0[98] = 16'b0000000000000000; P_DAT0[99] = 16'b0000000000000000;
	P_DAT0[100] = 16'b0000000000000000; P_DAT0[101] = 16'b0000000000000000; P_DAT0[102] = 16'b0000000000000000; P_DAT0[103] = 16'b0000000000000000;
	P_DAT0[104] = 16'b0000000000000000; P_DAT0[105] = 16'b0000000000000000; P_DAT0[106] = 16'b0000000000000000; P_DAT0[107] = 16'b0000000000000000;
	P_DAT0[108] = 16'b0000000000000000; P_DAT0[109] = 16'b0000000000000000; P_DAT0[110] = 16'b0000000000000000; P_DAT0[111] = 16'b0000000000000000;
	P_DAT0[112] = 16'b0000000000000000; P_DAT0[113] = 16'b0000000000000000; P_DAT0[114] = 16'b0000000000000000; P_DAT0[115] = 16'b0000000000000000;
	P_DAT0[116] = 16'b0000000000000000; P_DAT0[117] = 16'b0000000000000000; P_DAT0[118] = 16'b0000000000000000; P_DAT0[119] = 16'b0000000000000000;
	P_DAT0[120] = 16'b0000000000000000; P_DAT0[121] = 16'b0000000000000000; P_DAT0[122] = 16'b0000000000000000; P_DAT0[123] = 16'b0000000000000000;
	P_DAT0[124] = 16'b0000000000000000; P_DAT0[125] = 16'b0000000000000000; P_DAT0[126] = 16'b0000000000000000; P_DAT0[127] = 16'b0000000011111111;
	P_DAT0[128] = 16'b1100000000000000; P_DAT0[129] = 16'b0000000000000000; P_DAT0[130] = 16'b0000000000000000; P_DAT0[131] = 16'b0000000000000000;
	P_DAT0[132] = 16'b0000000000000000; P_DAT0[133] = 16'b0000000000000000; P_DAT0[134] = 16'b0000000000000000; P_DAT0[135] = 16'b0000000000000000;
	P_DAT0[136] = 16'b0000000000000000; P_DAT0[137] = 16'b0000000000000000; P_DAT0[138] = 16'b0000000000000000; P_DAT0[139] = 16'b0000000000000000;
	P_DAT0[140] = 16'b0000110000000000; P_DAT0[141] = 16'b0000110000000000; P_DAT0[142] = 16'b0000110000000000; P_DAT0[143] = 16'b0000110000000000;
	P_DAT0[144] = 16'b0001101110000000; P_DAT0[145] = 16'b0001101110000000; P_DAT0[146] = 16'b0001101110000000; P_DAT0[147] = 16'b0001101110000000;
	P_DAT0[148] = 16'b0000111110000000; P_DAT0[149] = 16'b0000111110000000; P_DAT0[150] = 16'b0000111110000000; P_DAT0[151] = 16'b0000111110000000;
	P_DAT0[152] = 16'b0000011100000000; P_DAT0[153] = 16'b0000011100000000; P_DAT0[154] = 16'b0000011100000000; P_DAT0[155] = 16'b0000011100000000;
	P_DAT0[156] = 16'b0000000000000000; P_DAT0[157] = 16'b0000000000000000; P_DAT0[158] = 16'b0000000000000000; P_DAT0[159] = 16'b0000000000000000;
	P_DAT0[160] = 16'b0000000000000000; P_DAT0[161] = 16'b0000000000000000; P_DAT0[162] = 16'b0000000000000000; P_DAT0[163] = 16'b0000000000000000;
	P_DAT0[164] = 16'b0000000000000000; P_DAT0[165] = 16'b0000000000000000; P_DAT0[166] = 16'b0001000000000000; P_DAT0[167] = 16'b0000000000000000;
	P_DAT0[168] = 16'b0000000000000000; P_DAT0[169] = 16'b0000000000000000; P_DAT0[170] = 16'b0000100000000000; P_DAT0[171] = 16'b0000000000000000;
	P_DAT0[172] = 16'b0000000000000000; P_DAT0[173] = 16'b0000000000000000; P_DAT0[174] = 16'b0000010000000000; P_DAT0[175] = 16'b0000000000000000;
	P_DAT0[176] = 16'b0000000000000000; P_DAT0[177] = 16'b0000000000000000; P_DAT0[178] = 16'b0000001000000000; P_DAT0[179] = 16'b0000000000000000;
	P_DAT0[180] = 16'b0000000000000000; P_DAT0[181] = 16'b0000000000000000; P_DAT0[182] = 16'b0000000000000000; P_DAT0[183] = 16'b0000000000000000;
	P_DAT0[184] = 16'b0000000000000000; P_DAT0[185] = 16'b0000000000000000; P_DAT0[186] = 16'b0000000000000000; P_DAT0[187] = 16'b0000000000000000;
	P_DAT0[188] = 16'b0000000000000000; P_DAT0[189] = 16'b0000000000000000; P_DAT0[190] = 16'b0000000000000000; P_DAT0[191] = 16'b0000000000000000;
	P_DAT0[192] = 16'b0000000000000000; P_DAT0[193] = 16'b0000000000000000; P_DAT0[194] = 16'b0000000000000000; P_DAT0[195] = 16'b0000000000000000;
	P_DAT0[196] = 16'b0000000000000000; P_DAT0[197] = 16'b0000000000000000; P_DAT0[198] = 16'b0000000000000000; P_DAT0[199] = 16'b0000000000000000;
	P_DAT0[200] = 16'b0000000000000000; P_DAT0[201] = 16'b0000000000000000; P_DAT0[202] = 16'b0000000000000000; P_DAT0[203] = 16'b0000000000000000;
	P_DAT0[204] = 16'b0000110000000000; P_DAT0[205] = 16'b0000111110000000; P_DAT0[206] = 16'b0000110000000000; P_DAT0[207] = 16'b0000110000000000;
	P_DAT0[208] = 16'b0001101110000000; P_DAT0[209] = 16'b0001101110000000; P_DAT0[210] = 16'b0001101110000000; P_DAT0[211] = 16'b0001101110000000;
	P_DAT0[212] = 16'b0000111110000000; P_DAT0[213] = 16'b0000111110000000; P_DAT0[214] = 16'b0000111110000000; P_DAT0[215] = 16'b0000111110000000;
	P_DAT0[216] = 16'b0000011100000000; P_DAT0[217] = 16'b0000011100000000; P_DAT0[218] = 16'b0000011100000000; P_DAT0[219] = 16'b0000011100000000;
	P_DAT0[220] = 16'b0000000000000000; P_DAT0[221] = 16'b0000000000000000; P_DAT0[222] = 16'b0000000000000000; P_DAT0[223] = 16'b0000000000000000;
	P_DAT0[224] = 16'b0000000000000000; P_DAT0[225] = 16'b0000000000000000; P_DAT0[226] = 16'b0000000000000000; P_DAT0[227] = 16'b0000000000000000;
	P_DAT0[228] = 16'b0000000000000000; P_DAT0[229] = 16'b0000000000000000; P_DAT0[230] = 16'b0000000000000000; P_DAT0[231] = 16'b0000000000000000;
	P_DAT0[232] = 16'b0000000000000000; P_DAT0[233] = 16'b0000000000000000; P_DAT0[234] = 16'b0000000000000000; P_DAT0[235] = 16'b0000000000000000;
	P_DAT0[236] = 16'b0000000000000000; P_DAT0[237] = 16'b0000000000000000; P_DAT0[238] = 16'b0000000000000000; P_DAT0[239] = 16'b0000000000000000;
	P_DAT0[240] = 16'b0000000000000000; P_DAT0[241] = 16'b0000000000000000; P_DAT0[242] = 16'b0000000000000000; P_DAT0[243] = 16'b0000000000000000;
	P_DAT0[244] = 16'b0000000000000000; P_DAT0[245] = 16'b0000000000000000; P_DAT0[246] = 16'b0000000000000000; P_DAT0[247] = 16'b0000000010000000;
	P_DAT0[248] = 16'b0000000000000000; P_DAT0[249] = 16'b0000000000000000; P_DAT0[250] = 16'b0000000000000000; P_DAT0[251] = 16'b0000000111000000;
	P_DAT0[252] = 16'b0000000000000000; P_DAT0[253] = 16'b0000000000000000; P_DAT0[254] = 16'b0000000000000000; P_DAT0[255] = 16'b0000000010000000;

	// Gosper's Glider Gun with eater
	P_DAT1[0] = 16'b0000000000000000; P_DAT1[1] = 16'b0000000000000000; P_DAT1[2] = 16'b0000000000000000; P_DAT1[3] = 16'b0000000000000000;
	P_DAT1[4] = 16'b0000000000000000; P_DAT1[5] =   16'b0000000001000000; P_DAT1[6] = 16'b0000000000000000; P_DAT1[7] = 16'b0000000000000000;
	P_DAT1[8] = 16'b0000000000000000; P_DAT1[9] =   16'b0000000101000000; P_DAT1[10] = 16'b0000000000000000; P_DAT1[11] = 16'b0000000000000000;
	P_DAT1[12] = 16'b0000000000000110; P_DAT1[13] = 16'b0000011000000000; P_DAT1[14] = 16'b0001100000000000; P_DAT1[15] = 16'b0000000000000000;
	P_DAT1[16] = 16'b0000000000001000; P_DAT1[17] = 16'b1000011000000000; P_DAT1[18] = 16'b0001100000000000; P_DAT1[19] = 16'b0000000000000000;
	P_DAT1[20] = 16'b0110000000010000; P_DAT1[21] = 16'b0100011000000000; P_DAT1[22] = 16'b0000000000000000; P_DAT1[23] = 16'b0000000000000000;
	P_DAT1[24] = 16'b0110000000010001; P_DAT1[25] = 16'b0110000101000000; P_DAT1[26] = 16'b0000000000000000; P_DAT1[27] = 16'b0000000000000000;
	P_DAT1[28] = 16'b0000000000010000; P_DAT1[29] = 16'b0100000001000000; P_DAT1[30] = 16'b0000000000000000; P_DAT1[31] = 16'b0000000000000000;
	P_DAT1[32] = 16'b0000000000001000; P_DAT1[33] = 16'b1000000000000000; P_DAT1[34] = 16'b0000000000000000; P_DAT1[35] = 16'b0000000000000000;
	P_DAT1[36] = 16'b0000000000000110; P_DAT1[37] = 16'b0000000000000000; P_DAT1[38] = 16'b0000000000000000; P_DAT1[39] = 16'b0000000000000000;
	P_DAT1[40] = 16'b0000000000000000; P_DAT1[41] = 16'b0000000000000000; P_DAT1[42] = 16'b0000000000000000; P_DAT1[43] = 16'b0000000000000000;
	P_DAT1[44] = 16'b0000000000000000; P_DAT1[45] = 16'b0000000000000000; P_DAT1[46] = 16'b0000000000000000; P_DAT1[47] = 16'b0000000000000000;
	P_DAT1[48] = 16'b0000000000000000; P_DAT1[49] = 16'b0000000000000000; P_DAT1[50] = 16'b0000000000000000; P_DAT1[51] = 16'b0000000000000000;
	P_DAT1[52] = 16'b0000000000000000; P_DAT1[53] = 16'b0000000000000000; P_DAT1[54] = 16'b0000000000000000; P_DAT1[55] = 16'b0000000000000000;
	P_DAT1[56] = 16'b0000000000000000; P_DAT1[57] = 16'b0000000000000000; P_DAT1[58] = 16'b0000000000000000; P_DAT1[59] = 16'b0000000000000000;
	P_DAT1[60] = 16'b0000000000000000; P_DAT1[61] = 16'b0000000000000000; P_DAT1[62] = 16'b0000000000000000; P_DAT1[63] = 16'b0000000000000000;
	P_DAT1[64] = 16'b0000000000000000; P_DAT1[65] = 16'b0000000000000000; P_DAT1[66] = 16'b0000000000000000; P_DAT1[67] = 16'b0000000000000000;
	P_DAT1[68] = 16'b0000000000000000; P_DAT1[69] = 16'b0000000000000000; P_DAT1[70] = 16'b0000000000000000; P_DAT1[71] = 16'b0000000000000000;
	P_DAT1[72] = 16'b0000000000000000; P_DAT1[73] = 16'b0000000000000000; P_DAT1[74] = 16'b0000000000000000; P_DAT1[75] = 16'b0000000000000000;
	P_DAT1[76] = 16'b0000000000000000; P_DAT1[77] = 16'b0000000000000000; P_DAT1[78] = 16'b0000000000000000; P_DAT1[79] = 16'b0000000000000000;
	P_DAT1[80] = 16'b0000000000000000; P_DAT1[81] = 16'b0000000000000000; P_DAT1[82] = 16'b0000000000000000; P_DAT1[83] = 16'b0000000000000000;
	P_DAT1[84] = 16'b0000000000000000; P_DAT1[85] = 16'b0000000000000000; P_DAT1[86] = 16'b0000000000000000; P_DAT1[87] = 16'b0000000000000000;
	P_DAT1[88] = 16'b0000000000000000; P_DAT1[89] = 16'b0000000000000000; P_DAT1[90] = 16'b0000000000000000; P_DAT1[91] = 16'b0000000000000000;
	P_DAT1[92] = 16'b0000000000000000; P_DAT1[93] = 16'b0000000000000000; P_DAT1[94] = 16'b0000000000000000; P_DAT1[95] = 16'b0000000000000000;
	P_DAT1[96] = 16'b0000000000000000; P_DAT1[97] = 16'b0000000000000000; P_DAT1[98] = 16'b0000000000000000; P_DAT1[99] = 16'b0000000000000000;
	P_DAT1[100] = 16'b0000000000000000; P_DAT1[101] = 16'b0000000000000000; P_DAT1[102] = 16'b0000000000000000; P_DAT1[103] = 16'b0000000000000000;
	P_DAT1[104] = 16'b0000000000000000; P_DAT1[105] = 16'b0000000000000000; P_DAT1[106] = 16'b0000000000000000; P_DAT1[107] = 16'b0000000000000000;
	P_DAT1[108] = 16'b0000000000000000; P_DAT1[109] = 16'b0000000000000000; P_DAT1[110] = 16'b0000000000000000; P_DAT1[111] = 16'b0000000000000000;
	P_DAT1[112] = 16'b0000000000000000; P_DAT1[113] = 16'b0000000000000000; P_DAT1[114] = 16'b0000000000000000; P_DAT1[115] = 16'b0000000000000000;
	P_DAT1[116] = 16'b0000000000000000; P_DAT1[117] = 16'b0000000000000000; P_DAT1[118] = 16'b0000000000000000; P_DAT1[119] = 16'b0000000000000000;
	P_DAT1[120] = 16'b0000000000000000; P_DAT1[121] = 16'b0000000000000000; P_DAT1[122] = 16'b0000110000000000; P_DAT1[123] = 16'b0000000000000000;
	P_DAT1[124] = 16'b0000000000000000; P_DAT1[125] = 16'b0000000000000000; P_DAT1[126] = 16'b0000110001000000; P_DAT1[127] = 16'b0000000000000000;
	P_DAT1[128] = 16'b0000000000000000; P_DAT1[129] = 16'b0000000000000000; P_DAT1[130] = 16'b0000000010100000; P_DAT1[131] = 16'b0000000000000000;
	P_DAT1[132] = 16'b0000000000000000; P_DAT1[133] = 16'b0000000000000000; P_DAT1[134] = 16'b0000000001010000; P_DAT1[135] = 16'b0000000000000000;
	P_DAT1[136] = 16'b0000000000000000; P_DAT1[137] = 16'b0000000000000000; P_DAT1[138] = 16'b0000000000010000; P_DAT1[139] = 16'b0000000000000000;
	P_DAT1[140] = 16'b0000000000000000; P_DAT1[141] = 16'b0000000000000000; P_DAT1[142] = 16'b0000000000011000; P_DAT1[143] = 16'b0000000000000000;
	P_DAT1[144] = 16'b0000000000000000; P_DAT1[145] = 16'b0000000000000000; P_DAT1[146] = 16'b0000000000000000; P_DAT1[147] = 16'b0000000000000000;
	P_DAT1[148] = 16'b0000000000000000; P_DAT1[149] = 16'b0000000000000000; P_DAT1[150] = 16'b0000000000000000; P_DAT1[151] = 16'b0000000000000000;
	P_DAT1[152] = 16'b0000000000000000; P_DAT1[153] = 16'b0000000000000000; P_DAT1[154] = 16'b0000000000000000; P_DAT1[155] = 16'b0000000000000000;
	P_DAT1[156] = 16'b0000000000000000; P_DAT1[157] = 16'b0000000000000000; P_DAT1[158] = 16'b0000000000000000; P_DAT1[159] = 16'b0000000000000000;
	P_DAT1[160] = 16'b0000000000000000; P_DAT1[161] = 16'b0000000000000000; P_DAT1[162] = 16'b0000000000000000; P_DAT1[163] = 16'b0000000000000000;
	P_DAT1[164] = 16'b0000000000000000; P_DAT1[165] = 16'b0000000000000000; P_DAT1[166] = 16'b0000000000000000; P_DAT1[167] = 16'b0000000000000000;
	P_DAT1[168] = 16'b0000000000000000; P_DAT1[169] = 16'b0000000000000000; P_DAT1[170] = 16'b0000000000000000; P_DAT1[171] = 16'b0000000000000000;
	P_DAT1[172] = 16'b0000000000000000; P_DAT1[173] = 16'b0000000000000000; P_DAT1[174] = 16'b0000000000000000; P_DAT1[175] = 16'b0000000000000000;
	P_DAT1[176] = 16'b0000000000000000; P_DAT1[177] = 16'b0000000000000000; P_DAT1[178] = 16'b0000000000000000; P_DAT1[179] = 16'b0000000000000000;
	P_DAT1[180] = 16'b0000000000000000; P_DAT1[181] = 16'b0000000000000000; P_DAT1[182] = 16'b0000000000000000; P_DAT1[183] = 16'b0000000000000000;
	P_DAT1[184] = 16'b0000000000000000; P_DAT1[185] = 16'b0000000000000000; P_DAT1[186] = 16'b0000000000000000; P_DAT1[187] = 16'b0000000000000000;
	P_DAT1[188] = 16'b0000000000000000; P_DAT1[189] = 16'b0000000000000000; P_DAT1[190] = 16'b0000000000000000; P_DAT1[191] = 16'b0000000000000000;
	P_DAT1[192] = 16'b0000000000000000; P_DAT1[193] = 16'b0000000000000000; P_DAT1[194] = 16'b0000000000000000; P_DAT1[195] = 16'b0000000000000000;
	P_DAT1[196] = 16'b0000000000000000; P_DAT1[197] = 16'b0000000000000000; P_DAT1[198] = 16'b0000000000000000; P_DAT1[199] = 16'b0000000000000000;
	P_DAT1[200] = 16'b0000000000000000; P_DAT1[201] = 16'b0000000000000000; P_DAT1[202] = 16'b0000000000000000; P_DAT1[203] = 16'b0000000000000000;
	P_DAT1[204] = 16'b0000000000000000; P_DAT1[205] = 16'b0000000000000000; P_DAT1[206] = 16'b0000000000000000; P_DAT1[207] = 16'b0000000000000000;
	P_DAT1[208] = 16'b0000000000000000; P_DAT1[209] = 16'b0000000000000000; P_DAT1[210] = 16'b0000000000000000; P_DAT1[211] = 16'b0000000000000000;
	P_DAT1[212] = 16'b0000000000000000; P_DAT1[213] = 16'b0000000000000000; P_DAT1[214] = 16'b0000000000000000; P_DAT1[215] = 16'b0000000000000000;
	P_DAT1[216] = 16'b0000000000000000; P_DAT1[217] = 16'b0000000000000000; P_DAT1[218] = 16'b0000000000000000; P_DAT1[219] = 16'b0000000000000000;
	P_DAT1[220] = 16'b0000000000000000; P_DAT1[221] = 16'b0000000000000000; P_DAT1[222] = 16'b0000000000000000; P_DAT1[223] = 16'b0000000000000000;
	P_DAT1[224] = 16'b0000000000000000; P_DAT1[225] = 16'b0000000000000000; P_DAT1[226] = 16'b0000000000000000; P_DAT1[227] = 16'b0000000000000000;
	P_DAT1[228] = 16'b0000000000000000; P_DAT1[229] = 16'b0000000000000000; P_DAT1[230] = 16'b0000000000000000; P_DAT1[231] = 16'b0000000000000000;
	P_DAT1[232] = 16'b0000000000000000; P_DAT1[233] = 16'b0000000000000000; P_DAT1[234] = 16'b0000000000000000; P_DAT1[235] = 16'b0000000000000000;
	P_DAT1[236] = 16'b0000000000000000; P_DAT1[237] = 16'b0000000000000000; P_DAT1[238] = 16'b0000000000000000; P_DAT1[239] = 16'b0000000000000000;
	P_DAT1[240] = 16'b0000000000000000; P_DAT1[241] = 16'b0000000000000000; P_DAT1[242] = 16'b0000000000000000; P_DAT1[243] = 16'b0000000000000000;
	P_DAT1[244] = 16'b0000000000000000; P_DAT1[245] = 16'b0000000000000000; P_DAT1[246] = 16'b0000000000000000; P_DAT1[247] = 16'b0000000000000000;
	P_DAT1[248] = 16'b0000000000000000; P_DAT1[249] = 16'b0000000000000000; P_DAT1[250] = 16'b0000000000000000; P_DAT1[251] = 16'b0000000000000000;
	P_DAT1[252] = 16'b0000000000000000; P_DAT1[253] = 16'b0000000000000000; P_DAT1[254] = 16'b0000000000000000; P_DAT1[255] = 16'b0000000000000000;

	// backrake
	P_DAT2[0] = 16'h0000; P_DAT2[1] = 16'h0000; P_DAT2[2] = 16'h0000; P_DAT2[3] = 16'h0000;
	P_DAT2[4] = 16'h0000; P_DAT2[5] =   16'h0000; P_DAT2[6] = 16'h0000; P_DAT2[7] = 16'h0000;
	P_DAT2[8] = 16'h0000; P_DAT2[9] =   16'h0000; P_DAT2[10] = 16'h0000; P_DAT2[11] = 16'h0000;
	P_DAT2[12] = 16'h0000; P_DAT2[13] = 16'h0000; P_DAT2[14] = 16'h0000; P_DAT2[15] = 16'h0000;
	P_DAT2[16] = 16'h0000; P_DAT2[17] = 16'h0000; P_DAT2[18] = 16'h0000; P_DAT2[19] = 16'h0000;
	P_DAT2[20] = 16'h0000; P_DAT2[21] = 16'h0000; P_DAT2[22] = 16'h0000; P_DAT2[23] = 16'h0000;
	P_DAT2[24] = 16'h0000; P_DAT2[25] = 16'h0000; P_DAT2[26] = 16'h0000; P_DAT2[27] = 16'h0000;
	P_DAT2[28] = 16'h0000; P_DAT2[29] = 16'h0000; P_DAT2[30] = 16'h0000; P_DAT2[31] = 16'h0000;
	P_DAT2[32] = 16'h0000; P_DAT2[33] = 16'h0000; P_DAT2[34] = 16'h0000; P_DAT2[35] = 16'h0000;
	P_DAT2[36] = 16'h0000; P_DAT2[37] = 16'h0000; P_DAT2[38] = 16'h0000; P_DAT2[39] = 16'h0000;
	P_DAT2[40] = 16'h0000; P_DAT2[41] = 16'h0000; P_DAT2[42] = 16'h0000; P_DAT2[43] = 16'h0000;
	P_DAT2[44] = 16'h0000; P_DAT2[45] = 16'h0000; P_DAT2[46] = 16'h0000; P_DAT2[47] = 16'h0000;
	P_DAT2[48] = 16'h0000; P_DAT2[49] = 16'h0000; P_DAT2[50] = 16'h0000; P_DAT2[51] = 16'h0000;
	P_DAT2[52] = 16'h0000; P_DAT2[53] = 16'h0000; P_DAT2[54] = 16'h0000; P_DAT2[55] = 16'h0000;
	P_DAT2[56] = 16'h0000; P_DAT2[57] = 16'h0000; P_DAT2[58] = 16'h0000; P_DAT2[59] = 16'h0000;
	P_DAT2[60] = 16'h0000; P_DAT2[61] = 16'h0000; P_DAT2[62] = 16'h0000; P_DAT2[63] = 16'h0000;
	P_DAT2[64] = 16'h0000; P_DAT2[65] = 16'h0000; P_DAT2[66] = 16'h0000; P_DAT2[67] = 16'h0000;
	P_DAT2[68] = 16'h0000; P_DAT2[69] = 16'h0000; P_DAT2[70] = 16'h0000; P_DAT2[71] = 16'h0000;
	P_DAT2[72] = 16'h0000; P_DAT2[73] = 16'h0000; P_DAT2[74] = 16'h0000; P_DAT2[75] = 16'h0000;
	P_DAT2[76] = 16'h0000; P_DAT2[77] = 16'h0000; P_DAT2[78] = 16'h0000; P_DAT2[79] = 16'h0000;
	P_DAT2[80] = 16'h0000; P_DAT2[81] = 16'h0000; P_DAT2[82] = 16'h0000; P_DAT2[83] = 16'h0000;
	P_DAT2[84] = 16'h0000; P_DAT2[85] = 16'h0000; P_DAT2[86] = 16'h0000; P_DAT2[87] = 16'h0000;
	P_DAT2[88] = 16'h0000; P_DAT2[89] = 16'h0000; P_DAT2[90] = 16'h0000; P_DAT2[91] = 16'h0000;
	P_DAT2[92] = 16'h0000; P_DAT2[93] = 16'h0000; P_DAT2[94] = 16'h0000; P_DAT2[95] = 16'h0000;
	P_DAT2[96] = 16'h0000; P_DAT2[97] = 16'h0000; P_DAT2[98] = 16'h0000; P_DAT2[99] = 16'h0000;
	P_DAT2[100] = 16'h0000; P_DAT2[101] = 16'b0000000111000000; P_DAT2[102] = 16'b0000011100000000; P_DAT2[103] = 16'h0000;
	P_DAT2[104] = 16'h0000; P_DAT2[105] = 16'b0000001000100000; P_DAT2[106] = 16'b0000100010000000; P_DAT2[107] = 16'h0000;
	P_DAT2[108] = 16'h0000; P_DAT2[109] = 16'b0000011000010000; P_DAT2[110] = 16'b0001000011000000; P_DAT2[111] = 16'h0000;
	P_DAT2[112] = 16'h0000; P_DAT2[113] = 16'b0000101011011000; P_DAT2[114] = 16'b0011011010100000; P_DAT2[115] = 16'h0000;
	P_DAT2[116] = 16'h0000; P_DAT2[117] = 16'b0001101000010110; P_DAT2[118] = 16'b1101000010110000; P_DAT2[119] = 16'h0000;
	P_DAT2[120] = 16'h0000; P_DAT2[121] = 16'b0010000100010010; P_DAT2[122] = 16'b1001000100001000; P_DAT2[123] = 16'h0000;
	P_DAT2[124] = 16'h0000; P_DAT2[125] = 16'b0000000000000010; P_DAT2[126] = 16'b1000000000000000; P_DAT2[127] = 16'h0000;
	P_DAT2[128] = 16'h0000; P_DAT2[129] = 16'b0011000000011010; P_DAT2[130] = 16'b1011000000011000; P_DAT2[131] = 16'h0000;
	P_DAT2[132] = 16'h0000; P_DAT2[133] = 16'b0000000000000010; P_DAT2[134] = 16'b1000000000000000; P_DAT2[135] = 16'h0000;
	P_DAT2[136] = 16'h0000; P_DAT2[137] = 16'b0000000011100000; P_DAT2[138] = 16'b0000111000000000; P_DAT2[139] = 16'h0000;
	P_DAT2[140] = 16'h0000; P_DAT2[141] = 16'b0000000010001000; P_DAT2[142] = 16'b0000001000000000; P_DAT2[143] = 16'h0000;
	P_DAT2[144] = 16'h0000; P_DAT2[145] = 16'b0000000010100001; P_DAT2[146] = 16'b1100000000000000; P_DAT2[147] = 16'h0000;
	P_DAT2[148] = 16'h0000; P_DAT2[149] = 16'b0000000000000010; P_DAT2[150] = 16'b0100001100000000; P_DAT2[151] = 16'h0000;
	P_DAT2[152] = 16'h0000; P_DAT2[153] = 16'b0000000000000000; P_DAT2[154] = 16'b0100000000000000; P_DAT2[155] = 16'h0000;
	P_DAT2[156] = 16'h0000; P_DAT2[157] = 16'b0000000000000100; P_DAT2[158] = 16'b0100000000000000; P_DAT2[159] = 16'h0000;
	P_DAT2[160] = 16'h0000; P_DAT2[161] = 16'b0000000000000100; P_DAT2[162] = 16'b0100000000000000; P_DAT2[163] = 16'h0000;
	P_DAT2[164] = 16'h0000; P_DAT2[165] = 16'b0000000000000000; P_DAT2[166] = 16'b0100000000000000; P_DAT2[167] = 16'h0000;
	P_DAT2[168] = 16'h0000; P_DAT2[169] = 16'b0000000000000010; P_DAT2[170] = 16'b1000000000000000; P_DAT2[171] = 16'h0000;
	P_DAT2[172] = 16'h0000; P_DAT2[173] = 16'h0000; P_DAT2[174] = 16'h0000; P_DAT2[175] = 16'h0000;
	P_DAT2[176] = 16'h0000; P_DAT2[177] = 16'h0000; P_DAT2[178] = 16'h0000; P_DAT2[179] = 16'h0000;
	P_DAT2[180] = 16'h0000; P_DAT2[181] = 16'h0000; P_DAT2[182] = 16'h0000; P_DAT2[183] = 16'h0000;
	P_DAT2[184] = 16'h0000; P_DAT2[185] = 16'h0000; P_DAT2[186] = 16'h0000; P_DAT2[187] = 16'h0000;
	P_DAT2[188] = 16'h0000; P_DAT2[189] = 16'h0000; P_DAT2[190] = 16'h0000; P_DAT2[191] = 16'h0000;
	P_DAT2[192] = 16'h0000; P_DAT2[193] = 16'h0000; P_DAT2[194] = 16'h0000; P_DAT2[195] = 16'h0000;
	P_DAT2[196] = 16'h0000; P_DAT2[197] = 16'h0000; P_DAT2[198] = 16'h0000; P_DAT2[199] = 16'h0000;
	P_DAT2[200] = 16'h0000; P_DAT2[201] = 16'h0000; P_DAT2[202] = 16'h0000; P_DAT2[203] = 16'h0000;
	P_DAT2[204] = 16'h0000; P_DAT2[205] = 16'h0000; P_DAT2[206] = 16'h0000; P_DAT2[207] = 16'h0000;
	P_DAT2[208] = 16'h0000; P_DAT2[209] = 16'h0000; P_DAT2[210] = 16'h0000; P_DAT2[211] = 16'h0000;
	P_DAT2[212] = 16'h0000; P_DAT2[213] = 16'h0000; P_DAT2[214] = 16'h0000; P_DAT2[215] = 16'h0000;
	P_DAT2[216] = 16'h0000; P_DAT2[217] = 16'h0000; P_DAT2[218] = 16'h0000; P_DAT2[219] = 16'h0000;
	P_DAT2[220] = 16'h0000; P_DAT2[221] = 16'h0000; P_DAT2[222] = 16'h0000; P_DAT2[223] = 16'h0000;
	P_DAT2[224] = 16'h0000; P_DAT2[225] = 16'h0000; P_DAT2[226] = 16'h0000; P_DAT2[227] = 16'h0000;
	P_DAT2[228] = 16'h0000; P_DAT2[229] = 16'h0000; P_DAT2[230] = 16'h0000; P_DAT2[231] = 16'h0000;
	P_DAT2[232] = 16'h0000; P_DAT2[233] = 16'h0000; P_DAT2[234] = 16'h0000; P_DAT2[235] = 16'h0000;
	P_DAT2[236] = 16'h0000; P_DAT2[237] = 16'h0000; P_DAT2[238] = 16'h0000; P_DAT2[239] = 16'h0000;
	P_DAT2[240] = 16'h0000; P_DAT2[241] = 16'h0000; P_DAT2[242] = 16'h0000; P_DAT2[243] = 16'h0000;
	P_DAT2[244] = 16'h0000; P_DAT2[245] = 16'h0000; P_DAT2[246] = 16'h0000; P_DAT2[247] = 16'h0000;
	P_DAT2[248] = 16'h0000; P_DAT2[249] = 16'h0000; P_DAT2[250] = 16'h0000; P_DAT2[251] = 16'h0000;
	P_DAT2[252] = 16'h0000; P_DAT2[253] = 16'h0000; P_DAT2[254] = 16'h0000; P_DAT2[255] = 16'h0000;

	// Traffic Circle
	P_DAT3[0] = 16'h0000; P_DAT3[1] = 16'h0000; P_DAT3[2] = 16'h0000; P_DAT3[3] = 16'h0000;
	P_DAT3[4] = 16'h0000; P_DAT3[5] =   16'h0000; P_DAT3[6] = 16'h0000; P_DAT3[7] = 16'h0000;
	P_DAT3[8] = 16'h0000; P_DAT3[9] =   16'h0000; P_DAT3[10] = 16'h0000; P_DAT3[11] = 16'h0000;
	P_DAT3[12] = 16'h0000; P_DAT3[13] = 16'h0000; P_DAT3[14] = 16'h0000; P_DAT3[15] = 16'h0000;
	P_DAT3[16] = 16'h0000; P_DAT3[17] = 16'h0000; P_DAT3[18] = 16'h0000; P_DAT3[19] = 16'h0000;
	P_DAT3[20] = 16'h0000; P_DAT3[21] = 16'h0000; P_DAT3[22] = 16'h0000; P_DAT3[23] = 16'h0000;
	P_DAT3[24] = 16'h0000; P_DAT3[25] = 16'h0000; P_DAT3[26] = 16'h0000; P_DAT3[27] = 16'h0000;
	P_DAT3[28] = 16'h0000; P_DAT3[29] = 16'h0000; P_DAT3[30] = 16'h0000; P_DAT3[31] = 16'h0000;
	P_DAT3[32] = 16'b0000000000000000; P_DAT3[33] = 16'b0000000000000110; P_DAT3[34] = 16'b0001100000000000; P_DAT3[35] = 16'b0000000000000000;
	P_DAT3[36] = 16'b0000000000000000; P_DAT3[37] = 16'b0000000000000101; P_DAT3[38] = 16'b0010100000000000; P_DAT3[39] = 16'b0000000000000000;
	P_DAT3[40] = 16'b0000000000000000; P_DAT3[41] = 16'b0000000000000001; P_DAT3[42] = 16'b0010000000000000; P_DAT3[43] = 16'b0000000000000000;
	P_DAT3[44] = 16'b0000000000000000; P_DAT3[45] = 16'b0000000000000011; P_DAT3[46] = 16'b0011000000000000; P_DAT3[47] = 16'b0000000000000000;
	P_DAT3[48] = 16'b0000000000000000; P_DAT3[49] = 16'b0000000000000111; P_DAT3[50] = 16'b0011100000000000; P_DAT3[51] = 16'b0000000000000000;
	P_DAT3[52] = 16'b0000000000000000; P_DAT3[53] = 16'b0000000000000001; P_DAT3[54] = 16'b0010000000000000; P_DAT3[55] = 16'b0000000000000000;
	P_DAT3[56] = 16'b0000000000000000; P_DAT3[57] = 16'b0000000000000000; P_DAT3[58] = 16'b0000000100000000; P_DAT3[59] = 16'b0000000000000000;
	P_DAT3[60] = 16'b0000000000000000; P_DAT3[61] = 16'b0000000000000000; P_DAT3[62] = 16'b0000001011000000; P_DAT3[63] = 16'b0000000000000000;
	P_DAT3[64] = 16'b0000000000000000; P_DAT3[65] = 16'b0000000000000000; P_DAT3[66] = 16'b0000000000100000; P_DAT3[67] = 16'b0000000000000000;
	P_DAT3[68] = 16'b0000000000000000; P_DAT3[69] = 16'b0000000000000000; P_DAT3[70] = 16'b0010001001010000; P_DAT3[71] = 16'b0000000000000000;
	P_DAT3[72] = 16'b0000000000000000; P_DAT3[73] = 16'b0000000000000000; P_DAT3[74] = 16'b0010000010010000; P_DAT3[75] = 16'b0000000000000000;
	P_DAT3[76] = 16'b0000000000000000; P_DAT3[77] = 16'b0000000000000000; P_DAT3[78] = 16'b0010000001100000; P_DAT3[79] = 16'b0000000000000000;
	P_DAT3[80] = 16'b0000000000000000; P_DAT3[81] = 16'b0110000000000000; P_DAT3[82] = 16'b0000000000000000; P_DAT3[83] = 16'b0000000000000000;
	P_DAT3[84] = 16'b0000000000000000; P_DAT3[85] = 16'b1001000000000011; P_DAT3[86] = 16'b1000111000000000; P_DAT3[87] = 16'b0000000000000000;
	P_DAT3[88] = 16'b0000000000000001; P_DAT3[89] = 16'b0101000000000000; P_DAT3[90] = 16'b0000000000000000; P_DAT3[91] = 16'b0000000000000000;
	P_DAT3[92] = 16'b0000000000000011; P_DAT3[93] = 16'b1010000000000000; P_DAT3[94] = 16'b0010000000000000; P_DAT3[95] = 16'b0000000000000000;
	P_DAT3[96] = 16'b0000000000000011; P_DAT3[97] = 16'b1000000000000000; P_DAT3[98] = 16'b0010000000000000; P_DAT3[99] = 16'b0000000000000000;
	P_DAT3[100] = 16'b0000000000000000; P_DAT3[101] = 16'b0000000000000000; P_DAT3[102] = 16'b0010000000000000; P_DAT3[103] = 16'b0000000000000000;
	P_DAT3[104] = 16'b0000000000000000; P_DAT3[105] = 16'b0000111000000000; P_DAT3[106] = 16'b0000000000000000; P_DAT3[107] = 16'b0000000000000000;
	P_DAT3[108] = 16'b0000000011001000; P_DAT3[109] = 16'b0000000000000111; P_DAT3[110] = 16'b0000000000000000; P_DAT3[111] = 16'b0000000000000000;
	P_DAT3[112] = 16'b0000000010011000; P_DAT3[113] = 16'b0010000010000000; P_DAT3[114] = 16'b0000000000000000; P_DAT3[115] = 16'b0000000000000000;
	P_DAT3[116] = 16'b0000000001111100; P_DAT3[117] = 16'b0010000010010000; P_DAT3[118] = 16'b0100000000000000; P_DAT3[119] = 16'b0001001100000000;
	P_DAT3[120] = 16'b0000000000000000; P_DAT3[121] = 16'b0010000010010000; P_DAT3[122] = 16'b0100000000000000; P_DAT3[123] = 16'b0001100100000000;
	P_DAT3[124] = 16'b0000000000000000; P_DAT3[125] = 16'b0000000000010000; P_DAT3[126] = 16'b0100000001110000; P_DAT3[127] = 16'b0011111000000000;
	P_DAT3[128] = 16'b0000000001111100; P_DAT3[129] = 16'b0000111000000000; P_DAT3[130] = 16'b0000000000000000; P_DAT3[131] = 16'b0000000000000000;
	P_DAT3[132] = 16'b0000000010011000; P_DAT3[133] = 16'b0000000000000111; P_DAT3[134] = 16'b0000000100000100; P_DAT3[135] = 16'b0000000000000000;
	P_DAT3[136] = 16'b0000000011001000; P_DAT3[137] = 16'b0000000000000000; P_DAT3[138] = 16'b0000000100000100; P_DAT3[139] = 16'b0011111000000000;
	P_DAT3[140] = 16'b0000000000000000; P_DAT3[141] = 16'b0000000000000000; P_DAT3[142] = 16'b0000000100000100; P_DAT3[143] = 16'b0001100100000000;
	P_DAT3[144] = 16'b0000000000000000; P_DAT3[145] = 16'b0000000000000000; P_DAT3[146] = 16'b0000000000000000; P_DAT3[147] = 16'b0001001100000000;
	P_DAT3[148] = 16'b0000000000000000; P_DAT3[149] = 16'b0000000000000000; P_DAT3[150] = 16'b0000000001110000; P_DAT3[151] = 16'b0000000000000000;
	P_DAT3[152] = 16'b0000000000000000; P_DAT3[153] = 16'b0000000000000000; P_DAT3[154] = 16'b0000000000000001; P_DAT3[155] = 16'b1000000000000000;
	P_DAT3[156] = 16'b0000000000000000; P_DAT3[157] = 16'b0000000000000000; P_DAT3[158] = 16'b0000000000000011; P_DAT3[159] = 16'b1000000000000000;
	P_DAT3[160] = 16'b0000000000000000; P_DAT3[161] = 16'b0000000000000000; P_DAT3[162] = 16'b0000000000000101; P_DAT3[163] = 16'b1000000000000000;
	P_DAT3[164] = 16'b0000000000000000; P_DAT3[165] = 16'b0000000000000000; P_DAT3[166] = 16'b0000000000001010; P_DAT3[167] = 16'b0000000000000000;
	P_DAT3[168] = 16'b0000000000000000; P_DAT3[169] = 16'b0000000000001110; P_DAT3[170] = 16'b0000000000001001; P_DAT3[171] = 16'b0000000000000000;
	P_DAT3[172] = 16'b0000000000000000; P_DAT3[173] = 16'b0000000000000000; P_DAT3[174] = 16'b0000000000000110; P_DAT3[175] = 16'b0000000000000000;
	P_DAT3[176] = 16'b0000000000000000; P_DAT3[177] = 16'b0000011000010010; P_DAT3[178] = 16'b0000000000000000; P_DAT3[179] = 16'b0000000000000000;
	P_DAT3[180] = 16'b0000000000000000; P_DAT3[181] = 16'b0000100100000000; P_DAT3[182] = 16'b0000000000000000; P_DAT3[183] = 16'b0000000000000000;
	P_DAT3[184] = 16'b0000000000000000; P_DAT3[185] = 16'b0000101010000000; P_DAT3[186] = 16'b0000000000000000; P_DAT3[187] = 16'b0000000000000000;
	P_DAT3[188] = 16'b0000000000000000; P_DAT3[189] = 16'b0000010010000000; P_DAT3[190] = 16'b0000000000000000; P_DAT3[191] = 16'b0000000000000000;
	P_DAT3[192] = 16'b0000000000000000; P_DAT3[193] = 16'b0000000001000000; P_DAT3[194] = 16'b0000000000000000; P_DAT3[195] = 16'b0000000000000000;
	P_DAT3[196] = 16'b0000000000000000; P_DAT3[197] = 16'b0000001010000000; P_DAT3[198] = 16'b0000000000000000; P_DAT3[199] = 16'b0000000000000000;
	P_DAT3[200] = 16'b0000000000000000; P_DAT3[201] = 16'b0000000000000100; P_DAT3[202] = 16'b1000000000000000; P_DAT3[203] = 16'b0000000000000000;
	P_DAT3[204] = 16'b0000000000000000; P_DAT3[205] = 16'b0000000000011100; P_DAT3[206] = 16'b1110000000000000; P_DAT3[207] = 16'b0000000000000000;
	P_DAT3[208] = 16'b0000000000000000; P_DAT3[209] = 16'b0000000000001100; P_DAT3[210] = 16'b1100000000000000; P_DAT3[211] = 16'b0000000000000000;
	P_DAT3[212] = 16'b0000000000000000; P_DAT3[213] = 16'b0000000000000100; P_DAT3[214] = 16'b1000000000000000; P_DAT3[215] = 16'b0000000000000000;
	P_DAT3[216] = 16'b0000000000000000; P_DAT3[217] = 16'b0000000000010100; P_DAT3[218] = 16'b1010000000000000; P_DAT3[219] = 16'b0000000000000000;
	P_DAT3[220] = 16'b0000000000000000; P_DAT3[221] = 16'b0000000000011000; P_DAT3[222] = 16'b0110000000000000; P_DAT3[223] = 16'b0000000000000000;
	P_DAT3[224] = 16'h0000; P_DAT3[225] = 16'h0000; P_DAT3[226] = 16'h0000; P_DAT3[227] = 16'h0000;
	P_DAT3[228] = 16'h0000; P_DAT3[229] = 16'h0000; P_DAT3[230] = 16'h0000; P_DAT3[231] = 16'h0000;
	P_DAT3[232] = 16'h0000; P_DAT3[233] = 16'h0000; P_DAT3[234] = 16'h0000; P_DAT3[235] = 16'h0000;
	P_DAT3[236] = 16'h0000; P_DAT3[237] = 16'h0000; P_DAT3[238] = 16'h0000; P_DAT3[239] = 16'h0000;
	P_DAT3[240] = 16'h0000; P_DAT3[241] = 16'h0000; P_DAT3[242] = 16'h0000; P_DAT3[243] = 16'h0000;
	P_DAT3[244] = 16'h0000; P_DAT3[245] = 16'h0000; P_DAT3[246] = 16'h0000; P_DAT3[247] = 16'h0000;
	P_DAT3[248] = 16'h0000; P_DAT3[249] = 16'h0000; P_DAT3[250] = 16'h0000; P_DAT3[251] = 16'h0000;
	P_DAT3[252] = 16'h0000; P_DAT3[253] = 16'h0000; P_DAT3[254] = 16'h0000; P_DAT3[255] = 16'h0000;

	// Achim's p144:
	P_DAT4[0] =  16'h0000; P_DAT4[1] =  16'h0000; P_DAT4[2] =  16'h0000; P_DAT4[3] =  16'h0000;
	P_DAT4[4] =  16'h0000; P_DAT4[5] =  16'h0000; P_DAT4[6] =  16'h0000; P_DAT4[7] =  16'h0000;
	P_DAT4[8] =  16'b0011000000000000; P_DAT4[9] =  16'b0000000000001100; P_DAT4[10] = 16'b0011000000000000; P_DAT4[11] = 16'b0000000000001100;
	P_DAT4[12] = 16'b0011000000000000; P_DAT4[13] = 16'b0000000000001100; P_DAT4[14] = 16'b0011000000000000; P_DAT4[15] = 16'b0000000000001100;
	P_DAT4[16] = 16'b0000000000000000; P_DAT4[17] = 16'b0000110000000000; P_DAT4[18] = 16'b0000000000110000; P_DAT4[19] = 16'b0000000000000000;
	P_DAT4[20] = 16'b0000000000000000; P_DAT4[21] = 16'b0001001000000000; P_DAT4[22] = 16'b0000000001001000; P_DAT4[23] = 16'b0000000000000000;
	P_DAT4[24] = 16'b0000000000000000; P_DAT4[25] = 16'b0000110000000000; P_DAT4[26] = 16'b0000000000110000; P_DAT4[27] = 16'b0000000000000000;
	P_DAT4[28] = 16'b0000000000000000; P_DAT4[29] = 16'b1000000000000000; P_DAT4[30] = 16'b0000000000000001; P_DAT4[31] = 16'b0000000000000000;
	P_DAT4[32] = 16'b0000000000000001; P_DAT4[33] = 16'b0100000000000000; P_DAT4[34] = 16'b0000000000000010; P_DAT4[35] = 16'b1000000000000000;
	P_DAT4[36] = 16'b0000000000000010; P_DAT4[37] = 16'b0010000000000000; P_DAT4[38] = 16'b0000000000000100; P_DAT4[39] = 16'b0100000000000000;
	P_DAT4[40] = 16'b0000000000000010; P_DAT4[41] = 16'b0100000000000000; P_DAT4[42] = 16'b0000000000000010; P_DAT4[43] = 16'b0100000000000000;
	P_DAT4[44] = 16'b0000000000000000; P_DAT4[45] = 16'b0000000000000000; P_DAT4[46] = 16'b0000000000000000; P_DAT4[47] = 16'b0000000000000000;
	P_DAT4[48] = 16'b0000000000000010; P_DAT4[49] = 16'b0100000000000000; P_DAT4[50] = 16'b0000000000000010; P_DAT4[51] = 16'b0100000000000000;
	P_DAT4[52] = 16'b0000000000000100; P_DAT4[53] = 16'b0100000000000000; P_DAT4[54] = 16'b0000000000000010; P_DAT4[55] = 16'b0010000000000000;
	P_DAT4[56] = 16'b0000000000000010; P_DAT4[57] = 16'b1000000000000000; P_DAT4[58] = 16'b0000000000000001; P_DAT4[59] = 16'b0100000000000000;
	P_DAT4[60] = 16'b0000000000000001; P_DAT4[61] = 16'b0000000000000000; P_DAT4[62] = 16'b0000000000000000; P_DAT4[63] = 16'b1000000000000000;
	P_DAT4[64] = 16'b0000000000110000; P_DAT4[65] = 16'b0000000000000000; P_DAT4[66] = 16'b0000000000000000; P_DAT4[67] = 16'b0000110000000000;
	P_DAT4[68] = 16'b0000000001001000; P_DAT4[69] = 16'b0000000000000000; P_DAT4[70] = 16'b0000000000000000; P_DAT4[71] = 16'b0001001000000000;
	P_DAT4[72] = 16'b0000000000110000; P_DAT4[73] = 16'b0000000000000000; P_DAT4[74] = 16'b0000000000000000; P_DAT4[75] = 16'b0000110000000000;
	P_DAT4[76] = 16'b0011000000000000; P_DAT4[77] = 16'b0000000000001100; P_DAT4[78] = 16'b0011000000000000; P_DAT4[79] = 16'b0000000000001100;
	P_DAT4[80] = 16'b0011000000000000; P_DAT4[81] = 16'b0000000000001100; P_DAT4[82] = 16'b0011000000000000; P_DAT4[83] = 16'b0000000000001100;
	P_DAT4[84] = 16'h0000; P_DAT4[85] = 16'h0000; P_DAT4[86] = 16'h0000; P_DAT4[87] = 16'h0000;
	P_DAT4[88] = 16'h0000; P_DAT4[89] = 16'h0000; P_DAT4[90] = 16'h0000; P_DAT4[91] = 16'h0000;
	P_DAT4[92] = 16'h0000; P_DAT4[93] = 16'h0000; P_DAT4[94] = 16'h0000; P_DAT4[95] = 16'h0000;
	P_DAT4[96] = 16'h0000; P_DAT4[97] = 16'h0000; P_DAT4[98] = 16'h0000; P_DAT4[99] = 16'h0000;
	P_DAT4[100] = 16'h0000; P_DAT4[101] = 16'h0000; P_DAT4[102] = 16'h0000; P_DAT4[103] = 16'h0000;
	P_DAT4[104] = 16'h0000; P_DAT4[105] = 16'h0000; P_DAT4[106] = 16'h0000; P_DAT4[107] = 16'h0000;
	P_DAT4[108] = 16'h0000; P_DAT4[109] = 16'h0000; P_DAT4[110] = 16'h0000; P_DAT4[111] = 16'h0000;
	P_DAT4[112] = 16'h0000; P_DAT4[113] = 16'h0000; P_DAT4[114] = 16'h0000; P_DAT4[115] = 16'h0000;
	P_DAT4[116] = 16'h0000; P_DAT4[117] = 16'h0000; P_DAT4[118] = 16'h0000; P_DAT4[119] = 16'h0000;
	P_DAT4[120] = 16'h0000; P_DAT4[121] = 16'h0000; P_DAT4[122] = 16'h0000; P_DAT4[123] = 16'h0000;
	P_DAT4[124] = 16'h0000; P_DAT4[125] = 16'h0000; P_DAT4[126] = 16'h0000; P_DAT4[127] = 16'h0000;
	P_DAT4[128] = 16'h0000; P_DAT4[129] = 16'h0000; P_DAT4[130] = 16'h0000; P_DAT4[131] = 16'h0000;
	P_DAT4[132] = 16'h0000; P_DAT4[133] = 16'h0000; P_DAT4[134] = 16'h0000; P_DAT4[135] = 16'h0000;
	P_DAT4[136] = 16'h0000; P_DAT4[137] = 16'h0000; P_DAT4[138] = 16'h0000; P_DAT4[139] = 16'h0000;
	P_DAT4[140] = 16'h0000; P_DAT4[141] = 16'h0000; P_DAT4[142] = 16'h0000; P_DAT4[143] = 16'h0000;
	P_DAT4[144] = 16'h0000; P_DAT4[145] = 16'h0000; P_DAT4[146] = 16'h0000; P_DAT4[147] = 16'h0000;
	P_DAT4[148] = 16'h0000; P_DAT4[149] = 16'h0000; P_DAT4[150] = 16'h0000; P_DAT4[151] = 16'h0000;
	P_DAT4[152] = 16'h0000; P_DAT4[153] = 16'h0000; P_DAT4[154] = 16'h0000; P_DAT4[155] = 16'h0000;
	P_DAT4[156] = 16'h0000; P_DAT4[157] = 16'h0000; P_DAT4[158] = 16'h0000; P_DAT4[159] = 16'h0000;
	P_DAT4[160] = 16'h0000; P_DAT4[161] = 16'h0000; P_DAT4[162] = 16'h0000; P_DAT4[163] = 16'h0000;
	P_DAT4[164] = 16'h0000; P_DAT4[165] = 16'h0000; P_DAT4[166] = 16'h0000; P_DAT4[167] = 16'h0000;
	P_DAT4[168] = 16'h0000; P_DAT4[169] = 16'h0000; P_DAT4[170] = 16'h0000; P_DAT4[171] = 16'h0000;
	P_DAT4[172] = 16'b0011000000000000; P_DAT4[173] = 16'b0000000000001100; P_DAT4[174] = 16'b0011000000000000; P_DAT4[175] = 16'b0000000000001100;
	P_DAT4[176] = 16'b0011000000000000; P_DAT4[177] = 16'b0000000000001100; P_DAT4[178] = 16'b0011000000000000; P_DAT4[179] = 16'b0000000000001100;
	P_DAT4[180] = 16'b0000000000110000; P_DAT4[181] = 16'b0000000000000000; P_DAT4[182] = 16'b0000000000000000; P_DAT4[183] = 16'b0000110000000000;
	P_DAT4[184] = 16'b0000000001001000; P_DAT4[185] = 16'b0000000000000000; P_DAT4[186] = 16'b0000000000000000; P_DAT4[187] = 16'b0001001000000000;
	P_DAT4[188] = 16'b0000000000110000; P_DAT4[189] = 16'b0000000000000000; P_DAT4[190] = 16'b0000000000000000; P_DAT4[191] = 16'b0000110000000000;
	P_DAT4[192] = 16'b0000000000000001; P_DAT4[193] = 16'b0000000000000000; P_DAT4[194] = 16'b0000000000000000; P_DAT4[195] = 16'b1000000000000000;
	P_DAT4[196] = 16'b0000000000000010; P_DAT4[197] = 16'b1000000000000000; P_DAT4[198] = 16'b0000000000000001; P_DAT4[199] = 16'b0100000000000000;
	P_DAT4[200] = 16'b0000000000000100; P_DAT4[201] = 16'b0100000000000000; P_DAT4[202] = 16'b0000000000000010; P_DAT4[203] = 16'b0010000000000000;
	P_DAT4[204] = 16'b0000000000000010; P_DAT4[205] = 16'b0100000000000000; P_DAT4[206] = 16'b0000000000000010; P_DAT4[207] = 16'b0100000000000000;
	P_DAT4[208] = 16'b0000000000000000; P_DAT4[209] = 16'b0000000000000000; P_DAT4[210] = 16'b0000000000000000; P_DAT4[211] = 16'b0000000000000000;
	P_DAT4[212] = 16'b0000000000000010; P_DAT4[213] = 16'b0100000000000000; P_DAT4[214] = 16'b0000000000000010; P_DAT4[215] = 16'b0100000000000000;
	P_DAT4[216] = 16'b0000000000000010; P_DAT4[217] = 16'b0010000000000000; P_DAT4[218] = 16'b0000000000000100; P_DAT4[219] = 16'b0100000000000000;
	P_DAT4[220] = 16'b0000000000000001; P_DAT4[221] = 16'b0100000000000000; P_DAT4[222] = 16'b0000000000000010; P_DAT4[223] = 16'b1000000000000000;
	P_DAT4[224] = 16'b0000000000000000; P_DAT4[225] = 16'b1000000000000000; P_DAT4[226] = 16'b0000000000000001; P_DAT4[227] = 16'b0000000000000000;
	P_DAT4[228] = 16'b0000000000000000; P_DAT4[229] = 16'b0000110000000000; P_DAT4[230] = 16'b0000000000110000; P_DAT4[231] = 16'b0000000000000000;
	P_DAT4[232] = 16'b0000000000000000; P_DAT4[233] = 16'b0001001000000000; P_DAT4[234] = 16'b0000000001001000; P_DAT4[235] = 16'b0000000000000000;
	P_DAT4[236] = 16'b0000000000000000; P_DAT4[237] = 16'b0000110000000000; P_DAT4[238] = 16'b0000000000110000; P_DAT4[239] = 16'b0000000000000000;
	P_DAT4[240] = 16'b0011000000000000; P_DAT4[241] = 16'b0000000000001100; P_DAT4[242] = 16'b0011000000000000; P_DAT4[243] = 16'b0000000000001100;
	P_DAT4[244] = 16'b0011000000000000; P_DAT4[245] = 16'b0000000000001100; P_DAT4[246] = 16'b0011000000000000; P_DAT4[247] = 16'b0000000000001100;
	P_DAT4[248] = 16'h0000; P_DAT4[249] = 16'h0000; P_DAT4[250] = 16'h0000; P_DAT4[251] = 16'h0000;
	P_DAT4[252] = 16'h0000; P_DAT4[253] = 16'h0000; P_DAT4[254] = 16'h0000; P_DAT4[255] = 16'h0000;

	// TODO: Add cool P_DAT 5 through 7

end

always @(posedge clk_24mhz)
begin
	if (state < 65 && state != 0)
	begin
		// Dont clock while latching and enabling
		CK <= ~CK;
	end

	half_div <= ~half_div;
	if (half_div) begin
		case (state)
			64:
			begin
				state <= state + 1;
				os_disp_addr <= 4*address + 0;
			end
			65:
			begin
				LA    <= 1;
				state <= state + 1;
				os_disp_addr <= 4*address + 1;

			end
			66:
			begin
				BL    <= 0;
				state <= state + 1;
				os_disp_addr <= 4*address + 2;
				r0_c0 <= os_t_data_out;
				r1_c0 <= os_b_data_out;
			end
			67:
			begin
				BL      <= 1;
				state   <= state + 1;
				os_disp_addr <= 4*address + 3;
				r0_c1 <= os_t_data_out;
				r1_c1 <= os_b_data_out;
			end
			68:
			begin
				{A4, A3, A2, A1, A0} <= address;
				CK                   <= 0;
				state                <= state + 1;
				LA                   <= 0;
				r0_c2 <= os_t_data_out;
				r1_c2 <= os_b_data_out;
			end
			69:
			begin
				r0_c3 <= os_t_data_out;
				r1_c3 <= os_b_data_out;
				state                <= state + 1;
			end
			70:
			begin
				address <= address + 1;
				state <= 0;
				// Arrange each 16 bits in the correct order or display nothing if the next
				// generation is not ready
				if (gol_state < 14) begin
					r0 <= 64'h0000000000000000;
					r1 <= 64'h0000000000000000;
				end else begin
					r0 <= {r0_c3[0], r0_c3[1], r0_c3[2], r0_c3[3], r0_c3[4], r0_c3[5], r0_c3[6], r0_c3[7], r0_c3[8], r0_c3[9], r0_c3[10], r0_c3[11], r0_c3[12], r0_c3[13], r0_c3[14], r0_c3[15],
						r0_c2[0], r0_c2[1], r0_c2[2], r0_c2[3], r0_c2[4], r0_c2[5], r0_c2[6], r0_c2[7], r0_c2[8], r0_c2[9], r0_c2[10], r0_c2[11], r0_c2[12], r0_c2[13], r0_c2[14], r0_c2[15],
						r0_c1[0], r0_c1[1], r0_c1[2], r0_c1[3], r0_c1[4], r0_c1[5], r0_c1[6], r0_c1[7], r0_c1[8], r0_c1[9], r0_c1[10], r0_c1[11], r0_c1[12], r0_c1[13], r0_c1[14], r0_c1[15],
						r0_c0[0], r0_c0[1], r0_c0[2], r0_c0[3], r0_c0[4], r0_c0[5], r0_c0[6], r0_c0[7], r0_c0[8], r0_c0[9], r0_c0[10], r0_c0[11], r0_c0[12], r0_c0[13], r0_c0[14], r0_c0[15]};
					r1 <= {r1_c3[0], r1_c3[1], r1_c3[2], r1_c3[3], r1_c3[4], r1_c3[5], r1_c3[6], r1_c3[7], r1_c3[8], r1_c3[9], r1_c3[10], r1_c3[11], r1_c3[12], r1_c3[13], r1_c3[14], r1_c3[15],
						r1_c2[0], r1_c2[1], r1_c2[2], r1_c2[3], r1_c2[4], r1_c2[5], r1_c2[6], r1_c2[7], r1_c2[8], r1_c2[9], r1_c2[10], r1_c2[11], r1_c2[12], r1_c2[13], r1_c2[14], r1_c2[15],
						r1_c1[0], r1_c1[1], r1_c1[2], r1_c1[3], r1_c1[4], r1_c1[5], r1_c1[6], r1_c1[7], r1_c1[8], r1_c1[9], r1_c1[10], r1_c1[11], r1_c1[12], r1_c1[13], r1_c1[14], r1_c1[15],
						r1_c0[0], r1_c0[1], r1_c0[2], r1_c0[3], r1_c0[4], r1_c0[5], r1_c0[6], r1_c0[7], r1_c0[8], r1_c0[9], r1_c0[10], r1_c0[11], r1_c0[12], r1_c0[13], r1_c0[14], r1_c0[15]};
				end
			end
			default:
			begin
				state     <= state + 1;
				R0        <= r0[horiz_cnt];
				R1        <= r1[horiz_cnt];
				G0        <= r0[horiz_cnt];
				G1        <= r1[horiz_cnt];
				B0        <= r0[horiz_cnt];
				B1        <= r1[horiz_cnt];
				horiz_cnt <= horiz_cnt + 1;
			end

		endcase
	end
end

endmodule
